module tb_chipmunks();

// Your testbench goes here.

endmodule: tb_chipmunks

// Any other simulation-only modules you need

